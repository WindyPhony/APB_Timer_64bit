module top(
	input wire sys_clk,
	input wire sys_rst_n,
	input wire tim_psel,
	input wire tim_pwrite,
	input wire tim_penable,
	input wire [11:0]tim_paddr,
	input wire [31:0]tim_pwdata,
	input wire dbg_mode,
	input wire [3:0] tim_pstrb,
	output wire [31:0]tim_prdata,
	output wire tim_pready,
	output wire tim_pslverr,
	output wire tim_int
);

wire WRITE_EN;
wire READ_EN;
wire div_en;
wire [3:0]div_val;
wire timer_en;
wire halt_ack;
wire err_div_val;
wire err_div_en;
wire cnt_en;
wire sel_wTDR0;
wire sel_wTDR1;
wire [31:0]DATA_TDR0;
wire [31:0]DATA_TDR1;
wire [63:0]COUNTER_VALUE;

register re(.CLK(sys_clk),
            .RST_N(sys_rst_n),
            .WRITE_EN(WRITE_EN),
            .READ_EN(READ_EN),
            .PADDR(tim_paddr),
            .PWDATA(tim_pwdata),
            .PSTRB(tim_pstrb),
            .COUNTER_VALUE(COUNTER_VALUE),
            .dbg_mode(dbg_mode),
            .halt_ack(halt_ack),
            .div_en(div_en),
            .div_val(div_val),
            .timer_en(timer_en),
            .sel_wTDR0(sel_wTDR0),
            .sel_wTDR1(sel_wTDR1),
            .PRDATA(tim_prdata),
            .PSLVERR(tim_pslverr),
            .tim_int(tim_int),
            .err_div_val_timer(err_div_val),
            .err_div_en(err_div_en),
            .DATA_TDR0(DATA_TDR0),	    
            .DATA_TDR1(DATA_TDR1),
	    .PREADY(tim_pready),
	    .PWRITE(tim_pwrite)	    
);

apb_slave as(.CLK(sys_clk),
	     .RST_N(sys_rst_n),
	     .PSEL(tim_psel),
	     .PENABLE(tim_penable),
	     .PWRITE(tim_pwrite),
	     .PREADY(tim_pready),
	     .WRITE_EN(WRITE_EN),
	     .READ_EN(READ_EN),
	     .PSLVERR(tim_pslverr)
);

counter_control cc(.CLK(sys_clk),
	           .RST_N(sys_rst_n),
		   .div_en(div_en),
		   .div_val(div_val),
		   .timer_en(timer_en),
	//	   .err_div_val(err_div_val),
	//	   .err_div_en(err_div_en),
		   .halt_ack(halt_ack),
		   .cnt_en(cnt_en)
);

counter co(.CLK(sys_clk),
	   .RST_N(sys_rst_n),
	   .sel_wTDR0(sel_wTDR0),
	   .sel_wTDR1(sel_wTDR1),
	   .timer_en(timer_en),
	   .cnt_en(cnt_en),
	   .DATA_TDR0(DATA_TDR0),
	   .DATA_TDR1(DATA_TDR1),
	   .COUNTER_VALUE(COUNTER_VALUE)
);
endmodule
