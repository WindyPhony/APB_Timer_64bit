module apb_slave (
	input wire CLK,
	input wire RST_N,
	input wire PSEL,
	input wire PENABLE,
	input wire PWRITE,
	input wire PSLVERR,
	output wire PREADY,
	output wire WRITE_EN,
	output wire READ_EN
);

reg ready;

always @(posedge CLK or negedge RST_N) begin
	if(!RST_N) begin
		ready <= 1'b0;
	end
	else begin
		ready <= PSEL & PENABLE & !ready;
	end
end

assign PREADY   = ready;
assign WRITE_EN = ready & (PWRITE & ~PSLVERR);
assign READ_EN  = ready & !PWRITE;

endmodule
